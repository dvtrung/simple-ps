module inp (
  input [15:0] inp,
  output [15:0] inpval
  );
  assign inpval = inp;
endmodule