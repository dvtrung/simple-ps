module hardware (
  input  clock,
  output led
  );
  
  assign led = clock;
endmodule
